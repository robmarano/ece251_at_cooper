module hello_tb;

  initial begin
  end // initial begin
endmodule